module moore_fsm_101 (input clk, input reset, input in, output reg out);     reg [1:0] state;     parameter S0 = 0, S1 = 1, S2 = 2;     always @(posedge clk) begin   if (reset) state <= S0;   else case (state)   S0: if (in) state <= S1;   S1: if (!in) state <= S2;   S2: if (in) state <= S1;   endcase   end     always @(state) begin   case (state)   S0: out = 0;   S1: out = 0;   S2: out = 1;   endcase   end     endmodule